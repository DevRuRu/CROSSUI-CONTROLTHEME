module biginteger

fn test_lshif