module biginteger

fn