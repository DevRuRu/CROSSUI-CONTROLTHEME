module biginteger

pub const (
	zero = BigIntege