module biginteger

fn test_lshift() {
	for a 