module bigin