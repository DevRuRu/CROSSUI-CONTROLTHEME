module biginteger

fn 