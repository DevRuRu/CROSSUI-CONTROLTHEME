module biginteger

fn test_multiply() {
	a := from_str('123456