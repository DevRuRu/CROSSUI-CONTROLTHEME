module biginteger

import strings

pub fn (big BigInteger) str() str