module biginteger

fn test_lshift() {
	for a in [i64(-777), 777] {
		a_big := from_i6