module biginteger

import math.bits

pub enum BigIntegerSign {
	negativ