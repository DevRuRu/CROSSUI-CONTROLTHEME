module bigint