module biginteger

pub fn