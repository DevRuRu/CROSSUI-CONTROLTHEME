module biginteger

fn test_divide_mod_big() {
	a := from_str('9876543123456789012345678