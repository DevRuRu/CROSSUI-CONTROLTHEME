module biginteger

pub fn (a BigI