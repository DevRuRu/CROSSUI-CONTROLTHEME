module biginteger

fn test_lshift() {
	for a in [i64(-777), 77