module biginteger

import strings

pub fn (big