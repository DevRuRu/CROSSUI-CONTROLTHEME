module biginteger

pub fn (a BigInteger) * (b BigInteger) BigInte