module bigintege