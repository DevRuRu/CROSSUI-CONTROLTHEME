module biginteger

fn test_from_str_neg_zero() {
