module biginteger

pub fn from_i8(i i8) BigInteger {
	return from_i64(