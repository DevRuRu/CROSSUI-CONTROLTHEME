module biginteger

im