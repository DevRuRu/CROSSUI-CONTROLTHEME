module biginteger

pub fn (big BigInteger) int() int {
	if big.sign ==