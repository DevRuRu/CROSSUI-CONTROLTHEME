module bi