module biginteger

pub fn (a BigInteger) * 