module biginteger

pub const (
	zero 