module biginteger

pub fn from