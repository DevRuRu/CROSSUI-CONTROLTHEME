module biginteger

fn test_multiply() {
	a := from_str('123456789012345678