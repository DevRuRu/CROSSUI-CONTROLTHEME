module biginteger

import ma