module biginteger

pub fn from_str(s