module biginteger

fn test_zero() {
	