module biginteger

pub fn from_str(str string) ?BigInteger {
	base := ten
	// V