module biginteger

pub