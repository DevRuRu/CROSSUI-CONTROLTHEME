module biginteger

pub const (
	zero = BigInteger{
		sign: .zero
		bits