module biginteger

pub con