module biginteger

pub fn (a BigInteger) * (b BigInte