module biginteger

pub fn (big BigIn