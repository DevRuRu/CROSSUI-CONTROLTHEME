
module biginteger

import math.bits

pub fn (a BigInteger) / (b BigInteger) BigInteger {