module biginteger

import strings

pu