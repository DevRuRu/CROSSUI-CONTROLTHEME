module biginteger

fn test_divide