module biginteger

pub 