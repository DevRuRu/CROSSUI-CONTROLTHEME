module biginteger

fn test_divide_mod_big() {
	a := from_str('98765