
module main

import os
import strconv
import hanabi1224.biginteger