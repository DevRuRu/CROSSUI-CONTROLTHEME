module biginteger

fn t