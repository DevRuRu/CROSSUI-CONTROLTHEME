module biginteger

fn test_divide_mod_big() {
	