module biginteger

fn test_divide_mod_big() {
	a := from_str('987654312345678901234567890') or { pa