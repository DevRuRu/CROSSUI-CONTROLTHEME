module biginteger

fn test_multiply