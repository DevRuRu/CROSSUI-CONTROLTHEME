module biginteger

pub fn (big BigInteger) int() 