module biginteger

import math.bits

pub enum Big