module biginteger