module biginteger
