module biginteger

pub fn from_str(str string) ?B