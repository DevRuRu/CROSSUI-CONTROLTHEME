
module biginteger
