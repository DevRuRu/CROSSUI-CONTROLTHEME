module biginteger

import strings

pub fn (big BigInteger) str() string {
	i