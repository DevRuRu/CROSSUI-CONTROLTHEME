module biginteger

p