module biginteger

import math.bits

pub e