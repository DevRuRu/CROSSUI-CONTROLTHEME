module biginteger

fn test