module biginteger

import math.bits

pub enum BigIntegerSign {
	negative = -1
	zero = 0
	positive =